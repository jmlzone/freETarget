module adc_drv(output logic sd, input pcm);

initial sd = 0;
int adrv, aint;
endmodule // adc_drv
